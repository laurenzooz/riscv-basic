module BLINKY (
  input CLK,
  input RESET,
  output [4:0] LEDS,
  input RXD, // emulates serial port
  output 02/08/2025

);


